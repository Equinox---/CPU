/*
 * Top Level Single-Cycle CPU module
 */


module SCMIPS(input sysclk,
				)