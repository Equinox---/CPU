//`timescale 1ns/1ps

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[30:2])
	0: data <= 32'b000010_00000000000000000000000011; // j Initial
	// illop:
	1: data <= 32'b000010_00000000000000000000010101; // j Interrupt
	// xadr:

	2: data <= 32'b000010_00000000000000000010100001; // j Exit1

	// Initial:
	3: data <= 32'b000000_00000_00000_01100_00000_100000; // add $t4 $0 $0
	4: data <= 32'b001111_00000_00100_0100000000000000; // lui $a0 0x4000
	5: data <= 32'b001000_00000_10000_0000000011111001; // addi $s0 $0 249
	6: data <= 32'b001000_00000_10001_0000000100100100; // addi $s1 $0 292
	7: data <= 32'b001000_00000_10010_0000001000110000; // addi $s2 $0 560
	8: data <= 32'b001000_00000_10011_0000010000011001; // addi $s3 $0 1049
	9: data <= 32'b001000_00000_11101_0000010000000000; // addi $sp $0 1024
	// Timer:

	24: data <= 32'b000011_00000000000000000010010110; // jal Normal
	25: data <= 32'b101011_00100_00000_0000000000001000; // sw $0 8($a0)
	26: data <= 32'b001111_00000_01000_1111111111111111; // lui $t0 0xffff
	27: data <= 32'b001001_01000_01000_1111111100000000; // addiu $t0 $t0 0xff00
	28: data <= 32'b101011_00100_01000_0000000000000000; // sw $t0 0($a0)
	29: data <= 32'b001001_01000_01000_0000000011111111; // addiu $t0 $t0 0xff
	30: data <= 32'b101011_00100_01000_0000000000000100; // sw $t0 4($a0)
	31: data <= 32'b001000_00000_01000_0000000000000011; // addi $t0 $0 3
	32: data <= 32'b101011_00100_01000_0000000000001000; // sw $t0 8($a0)
	33: data <= 32'b001000_00110_01101_0000000000000000; // addi $t5 $a2 0
	34: data <= 32'b001000_00111_01110_0000000000000000; // addi $t6 $a3 0
	35: data <= 32'b000000_01101_01110_01111_00000_100010; // sub $t7 $t5 $t6
	// Judge:
	36: data <= 32'b000100_01111_00000_0000000001110100; // beq $t7 $0 Exit
	37: data <= 32'b000001_01111_00000_0000000000000011; // bltz $t7 Negative
	// Positive:
	38: data <= 32'b000000_01110_00000_01101_00000_100000; // add $t5 $t6 $0
	39: data <= 32'b000000_01111_01110_01111_00000_100010; // sub $t7 $t7 $t6
	40: data <= 32'b000010_00000000000000000000100100; // j Judge
	// Negative:
	41: data <= 32'b000000_00000_01111_01110_00000_100010; // sub $t6 $0 $t7
	42: data <= 32'b000000_01101_01111_01111_00000_100000; // add $t7 $t5 $t7
	43: data <= 32'b000010_00000000000000000000100100; // j Judge
	// Interrupt:
	44: data <= 32'b100011_00100_01000_0000000000001000; // lw $t0 8($a0)
	45: data <= 32'b001100_01000_01000_1111111111111001; // andi $t0 $t0 0xfff9
	46: data <= 32'b101011_00100_01000_0000000000001000; // sw $t0 8($a0)
	47: data <= 32'b101011_11101_11111_0000000000000000; // sw $ra 0($sp)
	48: data <= 32'b000100_01100_00000_0000000000001110; // beq $t4 $0 First
	49: data <= 32'b001000_00000_01011_0000000000000001; // addi $t3 $0 1
	50: data <= 32'b000100_01100_01011_0000000000010010; // beq $t4 $t3 Second
	51: data <= 32'b001000_00000_01011_0000000000000010; // addi $t3 $0 2
	52: data <= 32'b000100_01100_01011_0000000000010110; // beq $t4 $t3 Third
	53: data <= 32'b001000_00000_01011_0000000000000011; // addi $t3 $0 3
	54: data <= 32'b000100_01100_01011_0000000000011010; // beq $t4 $t3 Fourth
	// Continue:
	55: data <= 32'b100011_11101_11111_0000000000000000; // lw $ra 0($sp)
	56: data <= 32'b101011_00100_00101_0000000000010100; // sw $a1 20($a0)
	57: data <= 32'b001001_00000_01001_0000000000000010; // addiu $t1 $0 2
	58: data <= 32'b100011_00100_01000_0000000000001000; // lw $t0 8($a0)
	59: data <= 32'b000000_01000_01001_01000_00000_100101; // or $t0 $t0 $t1
	60: data <= 32'b101011_00100_01000_0000000000001000; // sw $t0 8($a0)
	61: data <= 32'b001000_11010_11010_1111111111111100; // addi $26 $26 -4
	62: data <= 32'b000000_11010_00000_00000_00000_001000; // jr $26
	// First:
	63: data <= 32'b00000000000_00110_01000_11100_000000; // sll $t0 $a2 28
	64: data <= 32'b00000000000_01000_01000_11100_000010; // srl $t0 $t0 28
	65: data <= 32'b000011_00000000000000000001010111; // jal DigitalTube
	66: data <= 32'b001000_00101_00101_0000000010000000; // addi $a1 $a1 128
	67: data <= 32'b001000_00000_01100_0000000000000001; // addi $t4 $0 1
	68: data <= 32'b000010_00000000000000000000110111; // j Continue
	// Second:
	69: data <= 32'b00000000000_00110_01000_11000_000000; // sll $t0 $a2 24
	70: data <= 32'b00000000000_01000_01000_11100_000010; // srl $t0 $t0 28
	71: data <= 32'b000011_00000000000000000001010111; // jal DigitalTube
	72: data <= 32'b001000_00101_00101_0000000100000000; // addi $a1 $a1 256
	73: data <= 32'b001000_00000_01100_0000000000000010; // addi $t4 $0 2
	74: data <= 32'b000010_00000000000000000000110111; // j Continue
	// Third:
	75: data <= 32'b00000000000_00111_01000_11100_000000; // sll $t0 $a3 28
	76: data <= 32'b00000000000_01000_01000_11100_000010; // srl $t0 $t0 28
	77: data <= 32'b000011_00000000000000000001010111; // jal DigitalTube
	78: data <= 32'b001000_00101_00101_0000001000000000; // addi $a1 $a1 512
	79: data <= 32'b001000_00000_01100_0000000000000011; // addi $t4 $0 3
	80: data <= 32'b000010_00000000000000000000110111; // j Continue
	// Fourth:
	81: data <= 32'b00000000000_00111_01000_11000_000000; // sll $t0 $a3 24
	82: data <= 32'b00000000000_01000_01000_11100_000010; // srl $t0 $t0 28
	83: data <= 32'b000011_00000000000000000001010111; // jal DigitalTube
	84: data <= 32'b001000_00101_00101_0000010000000000; // addi $a1 $a1 1024
	85: data <= 32'b001000_00000_01100_0000000000000000; // addi $t4 $0 0
	86: data <= 32'b000010_00000000000000000000110111; // j Continue
	// DigitalTube:
	87: data <= 32'b001000_01000_01001_1111111111110001; // addi $t1 $t0 -15
	88: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Fifteen
	89: data <= 32'b001000_01000_01001_1111111111110010; // addi $t1 $t0 -14
	90: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Fourteen
	91: data <= 32'b001000_01000_01001_1111111111110011; // addi $t1 $t0 -13
	92: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Thirteen
	93: data <= 32'b001000_01000_01001_1111111111110100; // addi $t1 $t0 -12
	94: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Twelve
	95: data <= 32'b001000_01000_01001_1111111111110101; // addi $t1 $t0 -11
	96: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Eleven
	97: data <= 32'b001000_01000_01001_1111111111110110; // addi $t1 $t0 -10
	98: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Ten
	99: data <= 32'b001000_01000_01001_1111111111110111; // addi $t1 $t0 -9
	100: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Nine
	101: data <= 32'b001000_01000_01001_1111111111111000; // addi $t1 $t0 -8
	102: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Eight
	103: data <= 32'b001000_01000_01001_1111111111111001; // addi $t1 $t0 -7
	104: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Seven
	105: data <= 32'b001000_01000_01001_1111111111111010; // addi $t1 $t0 -6
	106: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Six
	107: data <= 32'b001000_01000_01001_1111111111111011; // addi $t1 $t0 -5
	108: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Five
	109: data <= 32'b001000_01000_01001_1111111111111100; // addi $t1 $t0 -4
	110: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Four
	111: data <= 32'b001000_01000_01001_1111111111111101; // addi $t1 $t0 -3
	112: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Three
	113: data <= 32'b001000_01000_01001_1111111111111110; // addi $t1 $t0 -2
	114: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 Two
	115: data <= 32'b001000_01000_01001_1111111111111111; // addi $t1 $t0 -1
	116: data <= 32'b000100_01001_00000_0000000000011101; // beq $t1 $0 One
	117: data <= 32'b000100_01000_00000_0000000000011110; // beq $t0 $0 Zero
	// Fifteen:
	118: data <= 32'b001000_00000_00101_0000000000001110; // addi $a1 $0 14
	119: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Fourteen:
	120: data <= 32'b001000_00000_00101_0000000000000110; // addi $a1 $0 6
	121: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Thirteen:
	122: data <= 32'b001000_00000_00101_0000000000100001; // addi $a1 $0 33
	123: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Twelve:
	124: data <= 32'b001000_00000_00101_0000000001000110; // addi $a1 $0 70
	125: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Eleven:
	126: data <= 32'b001000_00000_00101_0000000000000011; // addi $a1 $0 3
	127: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Ten:
	128: data <= 32'b001000_00000_00101_0000000000001000; // addi $a1 $0 8
	129: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Nine:
	130: data <= 32'b001000_00000_00101_0000000000010000; // addi $a1 $0 16
	131: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Eight:
	132: data <= 32'b001000_00000_00101_0000000000000000; // addi $a1 $0 0
	133: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Seven:
	134: data <= 32'b001000_00000_00101_0000000001111000; // addi $a1 $0 120
	135: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Six:
	136: data <= 32'b001000_00000_00101_0000000000000010; // addi $a1 $0 2
	137: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Five:
	138: data <= 32'b001000_00000_00101_0000000000010010; // addi $a1 $0 18
	139: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Four:
	140: data <= 32'b001000_00000_00101_0000000000011001; // addi $a1 $0 25
	141: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Three:
	142: data <= 32'b001000_00000_00101_0000000000110000; // addi $a1 $0 48
	143: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Two:
	144: data <= 32'b001000_00000_00101_0000000000100100; // addi $a1 $0 36
	145: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// One:
	146: data <= 32'b001000_00000_00101_0000000001111001; // addi $a1 $0 121
	147: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Zero:
	148: data <= 32'b001000_00000_00101_0000000001000000; // addi $a1 $0 64
	149: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Normal:
	150: data <= 32'b00000000000_11111_11111_00001_000000; // sll $ra $ra 1
	151: data <= 32'b00000000000_11111_11111_00001_000010; // srl $ra $ra 1
	152: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	// Exit:
	153: data <= 32'b000000_01110_00000_00010_00000_100000; // add $v0 $t6 $0
	154: data <= 32'b101011_00100_00010_0000000000001100; // sw $v0 12($a0)
	// UART_Send:
	155: data <= 32'b101011_00100_00010_0000000000011000; // sw $v0 24($a0)
	156: data <= 32'b100011_00100_01001_0000000000100000; // lw $t1 32($a0)
	157: data <= 32'b00000000000_01001_01001_00011_000010; // srl $t1 $t1 3
	158: data <= 32'b00000000000_01001_01001_00011_000000; // sll $t1 $t1 3
	159: data <= 32'b001001_01001_01001_0000000000000111; // addiu $t1 $t1 7
	160: data <= 32'b101011_00101_01001_0000000000100000; // sw $t1 32($a1)
>>>>>>> origin/master
	default: data <= 32'b0;//00010_00000000000000000000000011;
endcase
endmodule
