/*
 * scan mode displayer
 */




module DisplayTube(
					input Reset_n,
					input CLK,
					input [11:0] digit,
					output [27:0] display
					);



endmodule