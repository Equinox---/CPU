`timescale 1ns/1ps

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[6:2])
	// main:
	0: data <= 32'b000010_00000000000000000000000011; // j Normal
	// illop:
	1: data <= 32'b000010_00000000000000000000010011; // j Interrupt
	// xadr:
	2: data <= 32'b000010_00000000000000000000010011; // j Exit
	// Normal:
	3: data <= 32'b000011_00000000000000000000010000; // jal Enable_Int
	4: data <= 32'b001111_00000_00010_0100000000000000; // lui $v0 0x4000
	5: data <= 32'b001001_00010_00010_0000000000010000; // addiu $v0 $v0 0x10
	6: data <= 32'b100011_00010_00100_0000000000000000; // lw $a0 0($v0)
	7: data <= 32'b000000_00100_00100_00101_00000_100000; // add $a1 $a0 $a0
	8: data <= 32'b001000_00101_00110_1111111111111111; // addi $a2 $a1 -1
	9: data <= 32'b000000_00101_00110_00110_00000_100010; // sub $a2 $a1 $a2
	10: data <= 32'b000101_00110_00101_0000000000000001; // bne $a2 $a1 try
	11: data <= 32'b001000_00000_00110_0000000000000000; // addi $a2 $zero 0
	// try:
	12: data <= 32'b000000_00110_00101_00110_00000_100101; // or $a2 $a2 $a1
	13: data <= 32'b001000_00000_00101_0000000000000101; // addi $a1 $0 5
	14: data <= 32'b000100_00101_00110_1111111111111101; // beq $a1 $a2 try
	15: data <= 32'b000010_00000000000000000000010011; // j Exit
	// Enable_Int:
	16: data <= 32'b00000000000_11111_11111_00001_000000; // sll $ra $ra 1
	17: data <= 32'b00000000000_11111_11111_00001_000010; // srl $ra $ra 1
	18: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	default: data <= 32'b000010_00000000000000000000000011;
endcase
endmodule
