//`timescale 1ns/1ps

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[30:2])
	0: data <= 32'b000010_00000000000000000000000011; // j Initial
	// illop:
	1: data <= 32'b000010_00000000000000000000010101; // j Interrupt
	// xadr:
	2: data <= 32'b000010_00000000000000000000111101; // j Exit1
	// Initial:
	3: data <= 32'b000000_00000_00000_01100_00000_100000; // add $t4 $0 $0
	4: data <= 32'b001111_00000_00100_0100000000000000; // lui $a0 0x4000
	5: data <= 32'b001000_00000_10000_0000000011111001; // addi $s0 $0 249
	6: data <= 32'b001000_00000_10001_0000000100100100; // addi $s1 $0 292
	7: data <= 32'b001000_00000_10010_0000001000110000; // addi $s2 $0 560
	8: data <= 32'b001000_00000_10011_0000010000011001; // addi $s3 $0 1049
	9: data <= 32'b001000_00000_11101_0000010000000000; // addi $sp $0 1024
	// Timer:
	10: data <= 32'b000011_00000000000000000000111010; // jal Normal
	11: data <= 32'b101011_00100_00000_0000000000001000; // sw $0 8($a0)
	12: data <= 32'b001111_00000_01000_1111111111111111; // lui $t0 65535
	13: data <= 32'b001001_01000_01000_1111111100000000; // addiu $t0 $t0 65280
	14: data <= 32'b101011_00100_01000_0000000000000000; // sw $t0 0($a0)
	15: data <= 32'b001111_00000_01000_1111111111111111; // lui $t0 65535
	16: data <= 32'b001001_01000_01000_1111111111111111; // addiu $t0 $t0 65535
	17: data <= 32'b101011_00100_01000_0000000000000100; // sw $t0 4($a0)
	18: data <= 32'b001000_00000_01000_0000000000000011; // addi $t0 $0 3
	19: data <= 32'b101011_00100_01000_0000000000001000; // sw $t0 8($a0)
	20: data <= 32'b000010_00000000000000000000111101; // j Exit1
	// Interrupt:
	21: data <= 32'b101011_11101_11111_0000000000000000; // sw $ra 0($sp)
	22: data <= 32'b100011_11101_01100_1111111111111100; // lw $t4 -4($sp)
	23: data <= 32'b100011_00100_01000_0000000000001000; // lw $t0 8($a0)
	24: data <= 32'b001100_01000_01000_1111111111111001; // andi $t0 $t0 65529
	25: data <= 32'b101011_00100_01000_0000000000001000; // sw $t0 8($a0)
	26: data <= 32'b000100_01100_00000_0000000000001111; // beq $t4 $0 First
	27: data <= 32'b001000_00000_01011_0000000000000001; // addi $t3 $0 1
	28: data <= 32'b000100_01100_01011_0000000000010001; // beq $t4 $t3 Second
	29: data <= 32'b001000_00000_01011_0000000000000010; // addi $t3 $0 2
	30: data <= 32'b000100_01100_01011_0000000000010011; // beq $t4 $t3 Third
	31: data <= 32'b001000_00000_01011_0000000000000011; // addi $t3 $0 3
	32: data <= 32'b000100_01100_01011_0000000000010101; // beq $t4 $t3 Fourth
	// Continue:
	33: data <= 32'b101011_00100_00101_0000000000010100; // sw $a1 20($a0)
	34: data <= 32'b100011_00100_01000_0000000000001000; // lw $t0 8($a0)
	35: data <= 32'b001000_00000_00101_0000000000000010; // addi $a1 $0 2
	36: data <= 32'b000000_01000_00101_01000_00000_100101; // or $t0 $t0 $a1
	37: data <= 32'b101011_00100_01000_0000000000001000; // sw $t0 8($a0)
	38: data <= 32'b100011_11101_11111_0000000000000000; // lw $ra 0($sp)
	39: data <= 32'b101011_11101_01100_1111111111111100; // sw $t4 -4($sp)
	40: data <= 32'b001000_11010_11010_1111111111111100; // addi $26 $26 -4
	41: data <= 32'b000000_11010_00000_00000_00000_001000; // jr $26
	// First:
	42: data <= 32'b000000_00000_10000_00101_00000_100000; // add $a1 $0 $s0
	43: data <= 32'b001000_00000_01100_0000000000000001; // addi $t4 $0 1
	44: data <= 32'b101011_00100_01100_0000000000001100; // sw $t4 12($a0)
	45: data <= 32'b000010_00000000000000000000100001; // j Continue
	// Second:
	46: data <= 32'b000000_00000_10001_00101_00000_100000; // add $a1 $0 $s1
	47: data <= 32'b001000_00000_01100_0000000000000010; // addi $t4 $0 2
	48: data <= 32'b101011_00100_01100_0000000000001100; // sw $t4 12($a0)
	49: data <= 32'b000010_00000000000000000000100001; // j Continue
	// Third:
	50: data <= 32'b000000_00000_10010_00101_00000_100000; // add $a1 $0 $s2
	51: data <= 32'b001000_00000_01100_0000000000000011; // addi $t4 $0 3
	52: data <= 32'b101011_00100_01100_0000000000001100; // sw $t4 12($a0)
	53: data <= 32'b000010_00000000000000000000100001; // j Continue
	// Fourth:
	54: data <= 32'b000000_00000_10011_00101_00000_100000; // add $a1 $0 $s3
	55: data <= 32'b000000_00000_00000_01100_00000_100000; // add $t4 $0 $0
	56: data <= 32'b101011_00100_01100_0000000000001100; // sw $t4 12($a0)
	57: data <= 32'b000010_00000000000000000000100001; // j Continue
	// Normal:
	58: data <= 32'b000000_00000_11111_11111_00001_000000; // sll $ra $ra 1
	59: data <= 32'b000000_00000_11111_11111_00001_000010; // srl $ra $ra 1
	60: data <= 32'b000000_11111_00000_00000_00000_001000; // jr $ra
	default: data <= 32'b0;//00010_00000000000000000000000011;
endcase
endmodule
